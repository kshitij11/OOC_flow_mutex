
module test_gen (reset, clk, req0, req1, grant0, grant1);

input reset, clk, grant0, grant1;
output req0, req1;

endmodule
