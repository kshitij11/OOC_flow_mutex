
module mutex2 (req0, req1, grant0, grant1);

output grant0, grant1;
input req0, req1;

endmodule
